library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all; 

library grlib; 
use grlib.amba.all; 
use grlib.stdlib.all; 
use grlib.devices.all; 

library gaisler; 
use gaisler.misc.all; 

library UNISIM; 
use UNISIM.VComponents.all; 
 
entity AHB_bridge is 
  port( 
    -- Clock and Reset ----------------- 
    clkm   : in  std_logic; 
    rstn   : in  std_logic; 
    -- AHB Master records -------------- 
    ahbmi  : in  ahb_mst_in_type; 
    ahbmo  : out ahb_mst_out_type; 
    -- ARM Cortex-M0 AHB-Lite signals --     
    HADDR  : in  std_logic_vector (31 downto 0); -- AHB transaction address 
    HSIZE  : in  std_logic_vector (2 downto 0);  -- AHB size: byte, half-word or word 
    HTRANS : in  std_logic_vector (1 downto 0);  -- AHB transfer: non-sequential only 
    HWDATA : in  std_logic_vector (31 downto 0); -- AHB write-data 
    HWRITE : in  std_logic;                      -- AHB write control 
    HRDATA : out std_logic_vector (31 downto 0); -- AHB read-data 
    HREADY : out std_logic                       -- AHB stall signal 
  ); 
end; 
 
architecture structural of AHB_bridge is 
 
--declare a component for state_machine 
component state_machine is
  port (
    -- Clock and reset
    clkm    : in std_logic;
    rstn    : in std_logic;
    -- Wierd stuff
    dmai    : out ahb_dma_in_type;
    dmao    : in ahb_dma_out_type;
    -- ARM Cortext-M0 AHB-Lite signals
    HADDR   : in std_logic_vector (31 downto 0);
    HSIZE   : in std_logic_vector (2 downto 0);
    HTRANS  : in std_logic_vector (1 downto 0);
    HWRITE  : in std_logic;
    HREADY  : out std_logic
  );
end component;
   
--declare a component for ahbmst 
component ahbmst is
  port(
    -- Clock and reset
    clkm : in std_logic;
    rstn : in std_logic;
    -- AHB fun things
    dmai : in  ahb_dma_in_type;
    dmao : out ahb_dma_out_type;
    ahbo : out ahb_mst_out_type;
    ahbi : in ahb_mst_in_type
  );
end component;  
 
--declare a component for data_swapper
component data_swapper is 
  port (
    dmao    : in ahb_dma_out_type;
    -- ARM Cortex-M0 AHB-Lite Signals
    HRDATA  : out std_logic_vector (31 downto 0)
  );
end component;   
       
signal dmai : ahb_dma_in_type; 
signal dmao : ahb_dma_out_type; 
 
begin 
 
--instantiate state_machine component and make the connections 
init_state_machine : state_machine
  port map (clkm, rstn, dmai, dmao, HADDR, HSIZE, HTRANS, HWRITE, HREADY);
 
--instantiate the ahbmst component and make the connections   
init_ahbmst : ahbmst
  port  map (clkm, rstn, dmai, dmao, ahbmo, ahbmi);
 
--instantiate the data_swapper component and make the connections 
init_data_swapper : data_swapper
  port map (dmao, HRDATA);
 
end structural;